module FPUnit #(
    parameter width = 32
)  // 32-bits for ARMv3
(
    input                  CLK,          // Connect to CPU clock
    input                  RESET,        // Connect to the reset of the ARM processor.
    input                  FP_Start,     // Multi-cycle Enable. The control unit should assert this when FADD or FMUL instruction is detected.
    input                  FPUnitOp,     // Multi-cycle Operation. "0" for Single Float Addition, "1" for Single Float Multiplication. Generated by Control unit.
    input      [width-1:0] FP_Operand1,
    input      [width-1:0] FP_Operand2,
    output     [width-1:0] Result,
    output reg             FP_Busy       // Set immediately when FP_Start is set. Cleared when the Results become ready. This bit can be used to stall the processor while multi-cycle operations are on.
);

    localparam IDLE = 1'b0;
    localparam COMPUTING = 1'b1;

    reg state, n_state;
    reg Done;
    // state machine
    always @(posedge CLK or posedge RESET) begin
        if (RESET) state <= IDLE;
        else state <= n_state;
    end

    always @(*) begin
        case (state)
            IDLE: begin
                if (FP_Start) begin
                    n_state = COMPUTING;
                    FP_Busy = 1'b1;
                end 
                else begin
                    n_state = IDLE;
                    FP_Busy = 1'b0;
                end
            end
            COMPUTING: begin
                if (~Done) begin
                    n_state = COMPUTING;
                    FP_Busy = 1'b1;
                end 
                else begin
                    n_state = IDLE;
                    FP_Busy = 1'b0;
                end
            end
        endcase
    end

    // Multi-cycle 
    always @(posedge CLK or posedge RESET) begin : COMPUTING_PROCESS  // process which does the actual computation
        if (RESET) begin
            Done <= 0;
        end  
        else if (state == IDLE) begin // state: IDLE
            if (n_state == COMPUTING) begin
                Done <= 0;
            end
        end  
        else if (n_state == COMPUTING) begin // state: COMPUTING
            if (~FPUnitOp) begin  // Single Float Addition

            end  
            else begin  // Single Float Multiplication
                
            end
        end
    end



endmodule
