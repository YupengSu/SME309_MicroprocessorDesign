module ControlUnit(
    input [31:0] Instr,
    input [3:0] ALUFlags,
    input CLK,

    output MemtoReg,
    output MemWrite,
    output ALUSrc,
    output [1:0] ImmSrc,
    output RegWrite,
    output [2:0] RegSrc,
    output [1:0] ALUControl,	
    output PCSrc,
    output M_Start,
    output MCycleOp,
    output M_Write
    ); 
    
    wire [3:0] Cond;
    wire PSC, RegW, MemW, NoWrite;
    wire [1:0] FlagW;
    wire M_W;

    assign Cond=Instr[31:28];

    CondLogic CondLogic1(
        CLK,
        PCS,
        RegW,
        MemW,
        NoWrite,
        FlagW,
        Cond,
        ALUFlags,
        M_W,

        PCSrc,
        RegWrite,
        MemWrite,
        M_Write
    );

    Decoder Decoder1(
        Instr,

        PCS,
        RegW,
        MemW,
        MemtoReg,
        ALUSrc,
        ImmSrc,
        RegSrc,
        ALUControl,
        FlagW,
        NoWrite,
        M_Start,
        MCycleOp,
        M_W
    );
endmodule